/* Copyright(C) 2020 Cobac.Net All Rights Reserved. */
/* chapter: 第2章など表示回路を扱う各章    */
/* project: pattern, chardisp, dipslayなど */
/* outline: VGA用パラメータ                */

/* VGA(640×480)パラメータ */
localparam HPERIOD = 10'd800;
localparam HFRONT  = 10'd16;
localparam HWIDTH  = 10'd96;
localparam HBACK   = 10'd48;

localparam VPERIOD = 10'd525;
localparam VFRONT  = 10'd10;
localparam VWIDTH  = 10'd2;
localparam VBACK   = 10'd33;
